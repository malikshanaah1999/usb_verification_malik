

int num_of_bytes = 10;